/*
Author    				: 	Junhan Lv
Email Address         	:    1322069095@qq.com
Filename             	:    counter.v
Data                 	:    2023-11-9
Description           	:    counter for 60.
Modification History    	:
Data            Author       Version         Change Description
=======================================================
23/11/9        Junhan Lv    1.0              Original
*/

module key_filter (
    input  wire clk,
    input  wire rst_n,
    input  wire key_in  
);

always @(posedge clk or negedge rst_n) begin
    


end


    
endmodule

