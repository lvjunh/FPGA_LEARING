`timescale 1ns/1ns
module test(
input [31:0] bus,
input sel,
output check
);
//*************code***********//




//*************code***********//
endmodule